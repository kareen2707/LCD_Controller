-- Master_Controller submodule
-- Creation date: 12/12/2018
-- Last modification: 29/12/2018
-- Version: 2.0

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Master_Controller is
	port(
		Clk	:	in  std_logic;
		Reset_n	: 	in std_logic;
		
		--Configuration registers
		Address				: 	in unsigned(31 downto 0);
		DataLength			: 	in unsigned(31 downto 0);
		BurstCount			: 	in unsigned(2 downto 0);
		Start		 		:	in std_logic; -- Maybe we don't need it
		Currently_writing		:	in std_logic; 
		Reading	 			:	out std_logic;
		
		--Signals connected to FIFO
		
		FIFO_Almost_full		:	in std_logic;
		WrFIFO				: 	out std_logic;
		WrData				:	out std_logic_vector(31 downto 0);
		
		
		--Avalon Master Signals
		AM_WaitRequest			: 	in std_logic;
		AM_ReadDataValid 		:	in std_logic;
		AM_ReadData			:	in std_logic_vector(31 downto 0);
		AM_Address			: 	out std_logic_vector(31 downto 0);
		AM_Read 			:	out std_logic;
		AM_BurstCount 			:	out std_logic_vector(2 downto 0));
end entity Master_Controller;

architecture behavioural of Master_Controller is

-- State definition

type state is (Idle, WaitPermission, WaitFifo, WaitData, WriteData, AcqData );
signal CurrentState: state;

-- Auxiliar constants and signals 

constant burstsize		: integer := 4;
signal en_count 		: std_logic;
signal counter 			: integer range 0 to burstsize :=4; -- Counter used for AM_ReadDataValid	
Signal TmpAddress		: unsigned(31 downto 0);
Signal TmpLength		: unsigned (31 downto 0);
Signal TmpBurstCount	: unsigned (2 downto 0);

	
Begin
	WrFIFO <= '0';

	AM_process: Process (Clk, Reset_n)
	Begin

	if (Reset_n = '0') then
		WrFIFO <= '0';
		AM_Read <= '0';
		TmpAddress <= (others => '0');
		TmpBurstCount <= (others => '0');
		TmpLength <= (others => '0');
		WrData <= (others => '0');
		Reading <= '0';
		CurrentState <= Idle;
		
	elsif rising_edge(Clk) then
		
		case CurrentState is
			when Idle =>

				if Start = '1' then
				--if DataLength /= X"0000_0000" then	--Starting if length is higher than zero
					TmpAddress <= Address;
					TmpLength <= DataLength;
					TmpBurstCount <= BurstCount;
					CurrentState <= WaitPermission;
				end if;

			when WaitPermission =>
				if Currently_writing = '0' then
					CurrentState <= WaitFifo;
					AM_Address <= std_logic_vector(TmpAddress);
					AM_BurstCount <= std_logic_vector(TmpBurstCount);
				end if;

			when WaitFifo =>

				if FIFO_Almost_full = '0' then 
					CurrentState <= WaitData;
					WrFIFO <= '1';					--Notifying we want to write into the FIFO
					AM_Read <= '1';					--Initializing the reading process
					Reading <= '1';					--Notifying the SRAM module is been used by LCD Controller
				end if;
				
			when WaitData =>

				if AM_ReadDataValid = '1' then		--We have readed a new data from SRAM
					counter <= counter - 1;			--Counting the times that ReadDataValid is high
					WrData <= AM_ReadData;			--Each reading contains information of 2 pixels (each pixel = 16b)
					if counter = 0 then
						CurrentState <= AcqData;
					else
						counter <= 4;
						CurrentState <= WriteData;
					end if;						
				end if;
			
			when WriteData =>

				if AM_WaitRequest = '0' then
					CurrentState <= AcqData;
					AM_Read <= '0';
					WrFIFO <= '0';
				end if;

			when AcqData =>

				if AM_ReadDataValid = '0' then
					CurrentState <= WaitPermission;
					Reading <= '0';
					if TmpLength /= 1 then
						TmpAddress <= TmpAddress + 1;
						TmpLength <= TmpLength - 1;
					else
						TmpAddress <= Address;
						TmpLength <= DataLength;
					end if;
				end if;

			
		end case;	

	end if;

end process AM_process;
	
end ;